library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
entity UART_TX is
  generic (
    CLKS_PER_BIT : integer := 115    
    );
  port (
    i_Clk       : in  std_logic;
    i_TX_DV     : in  std_logic;
    i_TX_Byte   : in  std_logic_vector(7 downto 0);
    o_TX_Active : out std_logic;
    o_TX_Serial : out std_logic;
    o_TX_Done   : out std_logic
    );
end UART_TX;
 
 
architecture RTL of UART_TX is
 
  type t_SM_Main is (s_Idle, s_TX_Start_Bit, s_TX_Data_Bits,
                     s_TX_Stop_Bit, s_Cleanup, D);
  signal current_state, next_state : t_SM_Main := s_Idle;
 
  signal r_Clk_Count : integer range 0 to CLKS_PER_BIT-1 := 0;
  signal r_Bit_Index : integer range 0 to 7 := 0;  -- 8 Bits Total
  signal r_TX_Data   : std_logic_vector(7 downto 0) := (others => '0');
  signal r_TX_Done   : std_logic := '0';

begin
   
  p_UART_TX : process (i_Clk)
  begin
     
    if rising_edge(i_Clk) then
         
      case next_state is
 
        when s_Idle =>
          o_TX_Active <= '0';
          o_TX_Serial <= '1';         -- Drive Line High for Idle
          r_TX_Done   <= '0';
          r_Clk_Count <= 0;
          r_Bit_Index <= 0;
          
          if i_TX_DV = '1' then
            r_TX_Data <= i_TX_Byte;
            
            next_state <= s_TX_Start_Bit;
          else
            current_state <= s_Idle;
          end if;

        when s_TX_Start_Bit =>
          o_TX_Active <= '1';
          o_TX_Serial <= '0';
          current_state <= s_TX_Start_Bit;
          next_state <= D;
        
         when s_TX_Data_Bits =>
          o_TX_Serial <= r_TX_Data(r_Bit_Index);
          current_state <= s_TX_Data_Bits;
          next_state <= D;
    
         when s_TX_Stop_Bit =>
          o_TX_Serial <= '1';
          current_state <= s_TX_Stop_Bit;
          next_state <= D;

          when s_Cleanup =>
          o_TX_Active <= '0';
          r_TX_Done   <= '1';
          next_state   <= s_Idle;

         when D =>
         if r_Clk_Count < CLKS_PER_BIT-1 then
            r_Clk_Count <= r_Clk_Count + 1;
            next_state <= current_state;          
          else
            r_Clk_Count <= 0;
                case current_state is
                    when s_Idle => next_state <= s_TX_Start_Bit;
                    when s_TX_Start_Bit => next_state <= s_TX_Data_Bits;
                    when s_TX_Data_Bits => 
                                          -- Check if we have sent out all bits
                                             if r_Bit_Index < 7 then
                                               r_Bit_Index <= r_Bit_Index + 1;
                                               next_state  <= s_TX_Data_Bits;
                                             else
                                               r_Bit_Index <= 0;
                                               next_state   <= s_TX_Stop_Bit;
                                             end if;

                                           next_state <= s_TX_Stop_Bit;
                    
                    when s_TX_Stop_Bit => next_state <= s_Cleanup; 
                    when others => 
                           next_state <= s_Idle;
                end case;
            
          end if;

 
        when others =>
          next_state <= s_Idle;
 
      end case;
    end if;
  end process p_UART_TX;
 
  o_TX_Done <= r_TX_Done;
   
end RTL;
    